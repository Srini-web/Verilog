module notg (
  input wire a,
  output wire out
);

  assign out = ~a;

endmodule
